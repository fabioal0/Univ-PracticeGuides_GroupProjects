Library IEEE;
use IEEE.STD_Logic_1164.all;

entity simulacao
end simulacao;

architecture proc of simulacao is

signal s_xout, s_xin , s_reset, s_clk: STD_Logic;

end proc;
